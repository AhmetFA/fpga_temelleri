`include "uvm_macros.svh"
`include "uart_interface.sv"
import uvm_pkg::*;
module testbench;

    import test_list::*;
    //////////////////////////////////////////////////////////////////////////////
    // Declaration of Local Fields
    //////////////////////////////////////////////////////////////////////////////
    time clock_period = 10ns;
    bit clock;
    bit reset;

    //////////////////////////////////////////////////////////////////////////////
    //clock generation
    //////////////////////////////////////////////////////////////////////////////
    initial begin
        clock=0;
        forever #(clock_period/2) clock=~clock;
     end
    //////////////////////////////////////////////////////////////////////////////
    //reset Generation : change may required while generating reset for 
    //                   synchronous/Asynchronous or Active low/Active high
    //////////////////////////////////////////////////////////////////////////////
    initial begin
        reset = 1;  
        #(clock_period* 5) reset =0;
    end


    //////////////////////////////////////////////////////////////////////////////
    /*********************starting the execution uvm phases**********************/
    //////////////////////////////////////////////////////////////////////////////
    initial begin
        run_test();
      end


    //////////////////////////////////////////////////////////////////////////////
    //creatinng instance of interface, inorder to connect DUT and testcase
    //////////////////////////////////////////////////////////////////////////////
    uart_interface uart_intf(clock,reset);
  
    //////////////////////////////////////////////////////////////////////////////
    /*********************uart DUT Instantation **********************************/
    //////////////////////////////////////////////////////////////////////////////
    top dut (
        .clock(clock),
        .reset(reset),
        .sw(uart_intf.sw),
        .rx_din(uart_intf.rx_din),
        .tx_dout(uart_intf.tx_dout),
        .tx_active(uart_intf.tx_active),
        .rx_active(uart_intf.rx_active)
    );
    //////////////////////////////////////////////////////////////////////////////
    /**********Set the Interface instance Using Configuration Database***********/
    //////////////////////////////////////////////////////////////////////////////
    initial begin
        uvm_config_db#(virtual uart_interface)::set(uvm_root::get(),"*","vif",uart_intf);
    end
    
endmodule