`ifndef uart_transaction 
`define uart_transaction

class uart_transaction extends uvm_sequence_item;
  //////////////////////////////////////////////////////////////////////////////
  // Declaration of uart transaction fields
  //////////////////////////////////////////////////////////////////////////////
   rand bit [2:0] sw;
   rand bit [7:0] uart_stim_data;//data that is sent to dut
   logic [7:0]  uart_mon_data;//data that is received from dut
  //////////////////////////////////////////////////////////////////////////////
  //Declaration of Utility and Field macros,
  //////////////////////////////////////////////////////////////////////////////
  `uvm_object_utils_begin(uart_transaction)
    `uvm_field_int(sw,UVM_ALL_ON)
    `uvm_field_int(uart_stim_data,UVM_ALL_ON)
    `uvm_field_int(uart_mon_data,UVM_ALL_ON)
  `uvm_object_utils_end
   
  //////////////////////////////////////////////////////////////////////////////
  //Constructor
  //////////////////////////////////////////////////////////////////////////////
  function new(string name = "uart_transaction");
    super.new(name);
  endfunction
  //////////////////////////////////////////////////////////////////////////////
  // Declaration of Constraints
  //////////////////////////////////////////////////////////////////////////////

   
endclass


`endif


